
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Bandpass_filter is
	port (
		clk		: in std_logic;
		reset		: in std_logic;
		
		sink_data	: in std_logic_vector(31 downto 0);
		sink_error	: in std_logic_vector(1 downto 0);
		sink_valid	: in std_logic;

		source_data	: out std_logic_vector(31 downto 0);
		source_error	: out std_logic_vector(1 downto 0);
		source_valid	: out std_logic);
end entity;

architecture Bandpass_filter_arch of Bandpass_filter is

signal x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, 
x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32	:	signed (31 downto 0);
signal b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15, b16, b17,
b18, b19, b20, b21, b22, b23, b24, b25, b26, b27, b28, b29, b30, b31, b32	:  signed (31 downto 0);
signal p0, p1, p2, p3, p4, p5, p6, p7, p8, p9, p10, p11, p12, p13, p14, p15, p16, p17,
p18, p19, p20, p21, p22, p23, p24, p25, p26, p27, p28, p29, p30, p31, p32	:  signed (63 downto 0);
--signal x1, x2, x3, x4	:	signed (31 downto 0);
--signal b1, b2, b3, b4	:  signed (31 downto 0);
--signal p1, p2, p3, p4	:  signed (63 downto 0);
signal xSum	:	signed (68 downto 0);
signal f1, f2, f3, f4	:	unsigned (7 downto 0);


begin	
	b0 <= "11111000110110001111100110000001";--c = -0.055878460364900601 * 2^31  
	b1 <= "00000010010101100001011100111000";--c =  0.018252279579649325 * 2^31  
	b2 <= "00000011111000001010010100010101";--c =  0.030293116644193555 * 2^31  
	b3 <= "00000101101001001011111000100000";--c =  0.044090047370205721 * 2^31  
	b4 <= "00000110101100110101000110001111";--c =  0.052347368941352591 * 2^31  
	b5 <= "00000110010010001001100010101101";--c =  0.049090465773250158 * 2^31  
	b6 <= "00000100000101101100101111001101";--c =  0.031945681634075115 * 2^31  
	b7 <= "00000000011010111100010101011111";--c =  0.0032889094309224119 * 2^31 
	b8 <= "11111100001011010010100000001000";--c = -0.029871936946877897 * 2^31  
	b9 <= "11111000100101011010101011100001";--c = -0.057932510524848629 * 2^31  
	b10 <= "11110110110110100010010010001011";--c = -0.071467811703315717 * 2^31  
	b11 <= "11110111101010001100001100010001";--c = -0.065162293077486513 * 2^31  
	b12 <= "11111010111110011000101100010110";--c = -0.039259542603369169 * 2^31  
	b13 <= "11111111111101001110110110011001";--c = -0.00033788705256632134 * 2^31
	b14 <= "00000101001011111011001000001100";--c =  0.040518051195146849 * 2^31  
	b15 <= "00001001001000010101010011101001";--c =  0.07132970205248966 * 2^31   
	b16 <= "00001010100101110111010010110100";--m =  0.082747066407391018 * 2^31 
	b17 <= "00001001001000010101010011101001";--
	b18 <= "00000101001011111011001000001100";--
	b19 <= "11111111111101001110110110011001";--
	b20 <= "11111010111110011000101100010110";--
	b21 <= "11110111101010001100001100010001";--
	b22 <= "11110110110110100010010010001011";--
	b23 <= "11111000100101011010101011100001";--
	b24 <= "11111100001011010010100000001000";--
	b25 <= "00000000011010111100010101011111";--
	b26 <= "00000100000101101100101111001101";--
	b27 <= "00000110010010001001100010101101";--
	b28 <= "00000110101100110101000110001111";--
	b29 <= "00000101101001001011111000100000";--
	b30 <= "00000011111000001010010100010101";--
	b31 <= "00000010010101100001011100111000";--
	b32 <= "11111000110110001111100110000001";--
	
	
	process (clk, reset)
	begin
	if (reset = '1') then
		x0 <= "00000000000000000000000000000000";
		x1 <= "00000000000000000000000000000000";
		x2 <= "00000000000000000000000000000000";
		x3 <= "00000000000000000000000000000000";
		x4 <= "00000000000000000000000000000000";
		x5 <= "00000000000000000000000000000000";
		x6 <= "00000000000000000000000000000000";
		x7 <= "00000000000000000000000000000000";
		x8 <= "00000000000000000000000000000000";
		x9 <= "00000000000000000000000000000000";
		x10 <= "00000000000000000000000000000000";
		x11 <= "00000000000000000000000000000000";
		x12 <= "00000000000000000000000000000000";
		x13 <= "00000000000000000000000000000000";
		x14 <= "00000000000000000000000000000000";
		x15 <= "00000000000000000000000000000000";
		x16 <= "00000000000000000000000000000000";
		x17 <= "00000000000000000000000000000000";
		x18 <= "00000000000000000000000000000000";
		x19 <= "00000000000000000000000000000000";
		x20 <= "00000000000000000000000000000000";
		x21 <= "00000000000000000000000000000000";
		x22 <= "00000000000000000000000000000000";
		x23 <= "00000000000000000000000000000000";
		x24 <= "00000000000000000000000000000000";
		x25 <= "00000000000000000000000000000000";
		x26 <= "00000000000000000000000000000000";
		x27 <= "00000000000000000000000000000000";
		x28 <= "00000000000000000000000000000000";
		x29 <= "00000000000000000000000000000000";
		x30 <= "00000000000000000000000000000000";
		x31 <= "00000000000000000000000000000000";
		x32 <= "00000000000000000000000000000000";
        elsif (clk'event and clk = '1') then
            
		x32 <= x31;
        	x31 <= x30;
       		x30 <= x29;
		x29 <= x28;
        	x28 <= x27;
       		x27 <= x26;
		x26 <= x25;
        	x25 <= x24;
       		x24 <= x23;
		x23 <= x22;
        	x22 <= x21;
       		x21 <= x20;
		x20 <= x19;
        	x19 <= x18;
       		x18 <= x17;
		x17 <= x16;
        	x16 <= x15;
       		x15 <= x14;
		x14 <= x13;
        	x13 <= x12;
       		x12 <= x11;
		x11 <= x10;
        	x10 <= x9;
       		x9 <= x8;
		x8 <= x7;
        	x7 <= x6;
       		x6 <= x5;
		x5 <= x4;
        	x4 <= x3;
       		x3 <= x2;
       		x2 <= x1;
            	x1 <= x0;
            	x0 <= signed (sink_data);

            	p32 <= x32 * b32;
            	p31 <= x31 * b31;
            	p30 <= x30 * b30;
            	p29 <= x29 * b29;
            	p28 <= x28 * b28;
            	p27 <= x27 * b27;
            	p26 <= x26 * b26;
            	p25 <= x25 * b25;
            	p24 <= x24 * b24;
            	p23 <= x23 * b23;
            	p22 <= x22 * b22;
            	p21 <= x21 * b21;
		p20 <= x20 * b20;
            	p19 <= x19 * b19;
            	p18 <= x18 * b18;
            	p17 <= x17 * b17;
            	p16 <= x16 * b16;
            	p15 <= x15 * b15;
            	p14 <= x14 * b14;
            	p13 <= x13 * b13;
            	p12 <= x12 * b12;
            	p11 <= x11 * b11;
		p10 <= x10 * b10;
            	p9 <= x9 * b9;
            	p8 <= x8 * b8;
            	p7 <= x7 * b7;
            	p6 <= x6 * b6;
            	p5 <= x5 * b5;
            	p4 <= x4 * b4;
            	p3 <= x3 * b3;
            	p2 <= x2 * b2;
            	p1 <= x1 * b1;
            	p0 <= x0 * b0;

            	xSum <= resize(p1,xSum'length) + resize(p2,xSum'length) + resize(p3,xSum'length) + resize(p4,xSum'length) + resize(p5,xSum'length) + resize(p6,xSum'length) + resize(p7,xSum'length) + 
			resize(p8,xSum'length) + resize(p9,xSum'length) + resize(p10,xSum'length) + resize(p11,xSum'length) + resize(p12,xSum'length) + resize(p13,xSum'length) + resize(p14,xSum'length) + 
			resize(p15,xSum'length) + resize(p16,xSum'length) + resize(p17,xSum'length) + resize(p18,xSum'length) + resize(p19,xSum'length) + resize(p20,xSum'length) + resize(p21,xSum'length) + 
			resize(p22,xSum'length) + resize(p23,xSum'length) + resize(p24,xSum'length) + resize(p25,xSum'length) + resize(p26,xSum'length) + resize(p27,xSum'length) + resize(p28,xSum'length) + 
			resize(p29,xSum'length) + resize(p30,xSum'length) + resize(p31,xSum'length) + resize(p32,xSum'length);
            	source_data	<= std_logic_vector(xSum(61 downto 30));
        end if;
	end process;

	--source_data <= sink_data;

end architecture;